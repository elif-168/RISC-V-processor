// 3 tane mux lazım
//pcTarget add??


//module instantiations 